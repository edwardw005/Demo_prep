// Code your design here
`include "Top_level0.sv"
`include "ALU.sv"
`include "CTRL.sv"
`include "data_mem.sv"
`include "data_mem0.sv"
`include "InstROM.sv"
`include "LUT.sv"
`include "ProgCtrl.sv"
`include "RegFile.sv"
`include "Top_level.sv"
