// Code your testbench here
// or browse Examples
`include "fltflt_no_rnd_tb.sv"