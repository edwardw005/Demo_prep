// Code your testbench here
// or browse Examples
`include "flt2fix_tb.sv"