// Code your design here
`include "data_mem.sv"
`include "flt2fix0.sv"
`include "ALU.sv"
`include "CRTL.sv"
`include "InstROM.sv"
`include "LUT.sv"
`include "ProgCtrl.sv"
`include "RegFile.sv"
`include "flt2fix.sv"
