// Code your design here
`include "data_mem0.sv"
`include "Top_level0.sv"
`include "ALU.sv"
`include "CRTL.sv"
`include "data_mem.sv"
`include "InstROM.sv"
`include "LUT.sv"
`include "ProgCtrl.sv"
`include "RegFile.sv"
`include "Top_level.sv"

