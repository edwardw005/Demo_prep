// Code your design here
`include "data_mem.sv"
`include "data_mem0.sv"
`include "Top_level.sv"
`include "ALU.sv"
`include "CTRL.sv"
`include "InstROM.sv"
`include "ProgCtrl.sv"
`include "RegFile.sv"
`include "Top_level0.sv"
