// Code your design here
`include "data_mem.sv"
`include "fltflt_no_rnd.sv"
`include "ALU.sv"
`include "CRTL.sv"
`include "InstROM.sv"
`include "LUT.sv"
`include "ProgCtrl.sv"
`include "RegFile.sv"
`include "fltflt0_no_rnd.sv"

